`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:42:44 03/08/2022 
// Design Name: 
// Module Name:    MuxComp 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module MuxComp(
    input [4:0] R_FLAG,
    input [2:0] SEL_F,
    output S_FLAG
    );


endmodule
